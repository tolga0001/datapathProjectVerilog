module processor;
  reg [31:0] pc; // 32-bit program counter
  reg clk; // clock
  reg [7:0] datmem[0:31], mem[0:31]; // 32-size data and instruction memory (8 bit(1 byte) for each location)
  output reg [2:0] statusP; // 210 => nzv
  wire [31:0] 
    dataa, // Read data 1 output of Register File
    datab, // Read data 2 output of Register File
    out2,  // Output of mux with ALUSrc control - mult2
    out3,  // Output of mux with MemToReg control - mult3
    out4,  // Output of mux with (Branch & ALUZero) control - mult4
    out5,  // Output of mux with jalpc control - mult5
    sum,   // ALU result
    extad, // Output of sign-extend unit
    adder1out, // Output of adder which adds PC and 4 - add1
    adder2out, // Output of adder which adds PC+4 and 2 shifted sign-extend result - add2
    sextad; // Output of shift left 2 unit

  wire [5:0] inst31_26; // 31-26 bits of instruction
  wire [4:0] 
    inst25_21, // 25-21 bits of instruction
    inst20_16, // 20-16 bits of instruction
    inst15_11, // 15-11 bits of instruction
    out1;      // Write data input of Register File

  wire [15:0] inst15_0; // 15-0 bits of instruction

  wire [31:0] instruc, // current instruction
    dpack; // Read data output of memory (data read from memory)

  wire [2:0] gout; // Output of ALU control unit

  wire zout, // Zero output of ALU
    pcsrc, // Output of AND gate with Branch and ZeroOut inputs
    // Control signals
    regdest, alusrc, memtoreg, regwrite, memread, memwrite, branch, aluop1, aluop0, jalpc;

  // 32-size register file (32 bit(1 word) for each register)
  reg [31:0] registerfile[0:31];

  integer i;

  // datamemory connections
  always @(posedge clk) begin
    if (memwrite) begin
      // sum stores address, datab stores the value to be written
      datmem[sum[4:0]+3] <= datab[7:0];
      datmem[sum[4:0]+2] <= datab[15:8];
      datmem[sum[4:0]+1] <= datab[23:16];
      datmem[sum[4:0]] <= datab[31:24];
    end
  end

  // instruction memory
  // 4-byte instruction
  assign instruc = {mem[pc[4:0]], mem[pc[4:0]+1], mem[pc[4:0]+2], mem[pc[4:0]+3]};
  assign inst31_26 = instruc[31:26];
  assign inst25_21 = instruc[25:21];
  assign inst20_16 = instruc[20:16];
  assign inst15_11 = instruc[15:11];
  assign inst15_0 = instruc[15:0];

  // registers
  assign dataa = registerfile[inst25_21]; // Read register 1
  assign datab = registerfile[inst20_16]; // Read register 2

  always @(posedge clk) begin
    if (regwrite) begin
      registerfile[out1] <= out3; // Write data to register
    end
  end

  // read data from memory, sum stores address
  assign dpack = {datmem[sum[4:0]], datmem[sum[4:0]+1], datmem[sum[4:0]+2], datmem[sum[4:0]+3]};

  // multiplexers
  // mux with RegDst control
  mult2_to_1_5 mult1(out1, instruc[20:16], instruc[15:11], regdest);

  // mux with control balv_sig (for selecting 31. reg as destination) added by Tolga
  mul2_to_1_32 mult2();

  // mux with ALUSrc control
  mult2_to_1_32 mult3(out2, datab, extad, alusrc);

  // mux with MemToReg control
  mult2_to_1_32 mult4(out3, sum, dpack, memtoreg);

  // mux with (blezal && R[rs] <= 0)
  mul2_to_1_32 mult5(); // it will be implemented for blezal

  // mux with (Branch & ALUZero) control
  mult2_to_1_32 mult6(out4, adder1out, adder2out, pcsrc);

  // mux with (jalpc) control added by Tolga
  mul2_to_1_32 mult7(out5, out4, adder1out, jalpc);

  // mux with (balv) control added by Tolga
  mul2_to_1_32 mult8(); // it will be implemented for balv

  // mux with (Brv) control added by Tolga
  mul2_to_1_32 mult9(); // it will be implemented for brv

  // mux with select nandi // added by Tolga TODO: It will be implemented
  mul2_to_1_32 mul10(); // it will be added for selecting zeroextend nandi according to nandi signal

  // load pc
  always @(negedge clk) begin
    pc <= out4;
  end

  // alu, adder and control logic connections
  // ALU unit
  alu32 alu1(sum, dataa, out2, zout, gout, statusP);

  // adder which adds PC and 4
  adder add1(pc, 32'h4, adder1out);

  // adder which adds PC+4 and 2 shifted sign-extend result
  adder add2(adder1out, sextad, adder2out);

  // Control unit TODO: jalpc eklencek
  control cont(instruc[31:26], regdest, alusrc, memtoreg, regwrite, memread, memwrite, branch, aluop1, aluop0, jalpc);

  // Sign extend unit
  signext sext(instruc[15:0], extad);

  // ALU control unit
  alucont acont(aluop1, aluop0, instruc[3], instruc[2], instruc[1], instruc[0], gout);

  // Shift-left 2 unit
  shift shift2(sextad, extad);

  // AND gate
  assign pcsrc = (branch && zout) || jalpc; // added by Tolga

  // initialize datamemory, instruction memory and registers
  // read initial data from files given in hex
  initial begin
    $readmemh("initDm.dat", datmem); // read Data Memory
    $readmemh("initIM.dat", mem); // read Instruction Memory
    $readmemh("initReg.dat", registerfile); // read Register File

    for (i = 0; i < 32; i = i + 1) begin
      $display("Instruction Memory[%0d]= %h  ", i, mem[i], "Data Memory[%0d]= %h   ", i, datmem[i], "Register[%0d]= %h", i, registerfile[i]);
    end
  end

  initial begin
    pc = 0;
    #400 $finish;
  end

  initial begin
    clk = 0;
    // 40 time unit for each cycle
    forever #20 clk = ~clk;
  end

  initial begin
    $monitor($time, "PC %h", pc, "  SUM %h", sum, "   INST %h", instruc[31:0], "   REGISTER %h %h %h %h ", registerfile[4], registerfile[5], registerfile[6], registerfile[1]);
  end
endmodule
